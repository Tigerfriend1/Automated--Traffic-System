// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition"
// CREATED		"Fri Dec 09 11:19:24 2022"

module tff_XXX(
	clk,
	din,
	rst,
	dout
);


input wire	clk;
input wire	din;
input wire	rst;
output reg	dout;

wire	SYNTHESIZED_WIRE_0;





always@(posedge clk or negedge rst)
begin
if (!rst)
	begin
	dout <= 0;
	end
else
	dout <= dout ^ SYNTHESIZED_WIRE_0;
end


trigger	b2v_inst1(
	.Din(din),
	.CLK(clk),
	.rst_n(rst),
	.Dout(SYNTHESIZED_WIRE_0));


endmodule
